module flow_led(
input  sys_clk,
input  rst_n,
output led


);

endmodule